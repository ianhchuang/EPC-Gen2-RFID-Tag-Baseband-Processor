/*
	*	Clock/Reset Generator
	*
	*	CRG controls all clock and reset signal of all modules
	*
	*	Clock gating is applied to all modules for saving the power dissipation
	*
	*	The clock signal of each module vibrates in the lowest frequency for saving the power dissipation
	*
	*	The constraints of clock gating is specified in the file bb_proc.tcl
*/


`timescale 1us / 1ns


module crg
(
output clk_crc5,
output clk_crc16,
output clk_blf,
output clk_cp,
output clk_prng,
output reg clk_frm,
output clk_fm0,
output reg clk_mil,
output clk_mem,
output rst_n,
output reg rst_for_new_package,
output rst_crc16,
output reg start_working,
input clk_200K,					// 200 KHz input clock generated from multivibrator
input clk_dpie,					// delayed PIE code
input pie_code,
input rst,
input dr,
input [1:0]m,
input en_crc5,
input en_crc16,
input en_2nd_clk_cp,
input en_prng_idol,
input en_prng_act,
input en_tx,
input en_if,
input packet_complete_sync,
input en_crc16_for_rpy,
input reply_complete,
input rd_complete,
input bs_complete
);


wire clk_200K_n;
wire clk_blf_n;
wire rst_for_cpu_crc16;
wire en_crc16_rpy;				// compute a CRC-16 of the replying data
wire clk_crc16_1;
wire clk_crc16_2;
wire clk_dr0;
wire en_cp_1;
wire en_cp_2;
wire clk_cp_1;
wire clk_cp_2;
wire en_prng_idol_for_clk;
wire clk_prng_idol;
wire clk_blf_for_tx;
wire clk_blf_half_for_tx;
wire clk_blf_quar_for_tx;
wire clk_blf_eigh_for_tx;


reg en_crc5_d;
reg en_crc16_d;
reg en_crc16_for_rpy_d;
reg [1:0]reply_complete_d;
reg clk_dr1;
reg [2:0]cnt_dr0_p;
reg [2:0]cnt_dr0_n;
reg clk_dr0_p;
reg clk_dr0_n;
reg [1:0]dr_d;
reg term_cp_1;
reg [1:0]en_2nd_clk_cp_d;
reg en_prng_idol_d;
reg bs_complete_d;
reg clk_blf_half;	// clock signal in half of BLF
reg clk_blf_quar;	// clock signal in quarter of BLF
reg clk_blf_eigh;	// clock signal in one eighth of BLF
reg en_tx_d;
reg rd_complete_d;


// --- start working when clock generated by multivibrator is oscillating ---
always@(posedge clk_200K or negedge rst_n) begin
	if(~rst_n) start_working <= 1'b0;
	else start_working <= 1'b1;
end


// --- generate global low-active asynchronous reset ---
assign rst_n = ~rst;


// --- generate reset signal for a new package ---
always@(negedge clk_dpie or negedge rst_n) begin
	if(~rst_n) rst_for_new_package <= 1'b1;
	else begin
		if(~pie_code) rst_for_new_package <= 1'b0;
		else rst_for_new_package <= 1'b1;
	end
end


// --- generate reset signal for CRC-16 ---
assign rst_for_cpu_crc16 = en_crc16_for_rpy & ~en_crc16_for_rpy_d;

assign rst_crc16 = rst_for_new_package & ~rst_for_cpu_crc16;


// --- generate clock signal of CRC-5 ---
always@(negedge clk_dpie or negedge rst_n) begin
	if(~rst_n) en_crc5_d <= 1'b0;
	else en_crc5_d <= en_crc5;
end

assign clk_crc5 = en_crc5_d & clk_dpie;


// --- generate clock signal of CRC-16 ---
always@(posedge clk_dpie or negedge rst_n) begin
	if(~rst_n) en_crc16_d <= 1'b0;
	else en_crc16_d <= en_crc16;
end

always@(negedge clk_frm or negedge rst_n) begin
	if(~rst_n) en_crc16_for_rpy_d <= 1'b0;
	else en_crc16_for_rpy_d <= en_crc16_for_rpy;
end

always@(negedge clk_frm or negedge rst_n) begin
	if(~rst_n) reply_complete_d <= 2'b0;
	else reply_complete_d <= {reply_complete_d[0], reply_complete};
end

assign en_crc16_rpy = en_crc16_for_rpy_d & ~reply_complete_d[1];

assign clk_crc16_1 = en_crc16_d & clk_dpie;

assign clk_crc16_2 = en_crc16_rpy & clk_frm;

assign clk_crc16 = en_crc16_for_rpy? clk_crc16_2 : clk_crc16_1;


// --- generate 100 KHz clock for DR = 1 (divide 2) ---
always@(posedge clk_200K or negedge rst_n) begin
	if(~rst_n) clk_dr1 <= 1'b0;
	else begin
		if(dr_d[1]) clk_dr1 <= ~clk_dr1;
	end
end


// --- generate 40 KHz clock for DR = 0 (divide 5) ---
assign clk_dr0 = clk_dr0_p | clk_dr0_n;

always@(posedge clk_200K or negedge rst_n) begin
	if(~rst_n) cnt_dr0_p <= 3'b0;
	else begin
		if(~dr_d[1]) begin
			if(cnt_dr0_p == 3'b100) cnt_dr0_p <= 3'b0;
			else cnt_dr0_p <= cnt_dr0_p + 3'b1;
		end
	end
end

assign clk_200K_n = ~clk_200K;

always@(posedge clk_200K_n or negedge rst_n) begin
	if(~rst_n) cnt_dr0_n <= 3'b0;
	else begin
		if(~dr_d[1]) begin
			if(cnt_dr0_n == 3'b100) cnt_dr0_n <= 3'b0;
			else cnt_dr0_n <= cnt_dr0_n + 3'b1;
		end
	end
end

always@(posedge clk_200K or negedge rst_n) begin
	if(~rst_n) clk_dr0_p <= 1'b0;
	else begin
		if(~dr_d[1]) begin
			if(cnt_dr0_p < 3'b010) clk_dr0_p <= 1'b1;
			else clk_dr0_p <= 1'b0;
		end
	end
end

always@(posedge clk_200K_n or negedge rst_n) begin
	if(~rst_n) clk_dr0_n <= 1'b0;
	else begin
		if(~dr_d[1]) begin
			if(cnt_dr0_n < 3'b010) clk_dr0_n <= 1'b1;
			else clk_dr0_n <= 1'b0;
		end
	end
end


// --- determine backscatter link frequency of clock ---
always@(posedge clk_blf or negedge rst_n) begin
	if(~rst_n) dr_d <= 0;
	else dr_d <= {dr_d[0], dr};
end

assign clk_blf = dr_d[1]? clk_dr1 : clk_dr0;


// --- generate clock signal of Command Processor ---
assign clk_blf_n = ~clk_blf;

always@(posedge clk_blf_n or negedge rst_n) begin
	if(~rst_n) term_cp_1 <= 1'b0;
	else term_cp_1 <= packet_complete_sync;
end

assign en_cp_1 = packet_complete_sync & ~term_cp_1;

always@(posedge clk_blf_n or negedge rst_n) begin
	if(~rst_n) en_2nd_clk_cp_d <= 2'b0;
	else en_2nd_clk_cp_d <= {en_2nd_clk_cp_d[0], en_2nd_clk_cp};
end

assign en_cp_2 = ~en_2nd_clk_cp_d[1] & en_2nd_clk_cp_d[0];

assign clk_cp_1 = clk_blf & en_cp_1;

assign clk_cp_2 = clk_blf & en_cp_2;

assign clk_cp = clk_cp_1 | clk_cp_2;


// --- generate clock signal of PRNG ---
always@(posedge clk_blf_n or negedge rst_n) begin
	if(~rst_n) en_prng_idol_d <= 1'b0;
	else en_prng_idol_d <= en_prng_idol;
end

assign clk_prng_idol = clk_blf & en_prng_idol_d;

assign clk_prng = start_working & (clk_prng_idol | en_prng_act);


// --- generate clock signal of Frame Generator ---
always@(posedge clk_blf_n or negedge rst_n) begin
	if(~rst_n) bs_complete_d <= 1'b0;
	else bs_complete_d <= bs_complete;
end

always@(posedge clk_blf or negedge rst_n) begin
	if(~rst_n) en_tx_d <= 1'b0;
	else en_tx_d <= en_tx;
end

always@(posedge clk_blf or negedge rst_n) begin
	if(~rst_n) clk_blf_half <= 1'b0;
	else if(en_tx & (m == 2'b01 | m == 2'b10 | m == 2'b11)) clk_blf_half <= ~clk_blf_half;
end

always@(posedge clk_blf_half or negedge rst_n) begin
	if(~rst_n) clk_blf_quar <= 1'b0;
	else if(en_tx & (m == 2'b10 | m == 2'b11)) clk_blf_quar <= ~clk_blf_quar;
end

always@(posedge clk_blf_quar or negedge rst_n) begin
	if(~rst_n) clk_blf_eigh <= 1'b0;
	else if(en_tx & m == 2'b11) clk_blf_eigh <= ~clk_blf_eigh;
end

assign clk_blf_for_tx = clk_blf & en_tx_d & ~bs_complete_d;

assign clk_blf_half_for_tx = clk_blf_half & ~bs_complete_d;

assign clk_blf_quar_for_tx = clk_blf_quar & ~bs_complete_d;

assign clk_blf_eigh_for_tx = clk_blf_eigh & ~bs_complete_d;

always@(*) begin
	if(en_tx) begin
		case(m)
			2'b00 : clk_frm = clk_blf_for_tx;
			2'b01 : clk_frm = clk_blf_half_for_tx;
			2'b10 : clk_frm = clk_blf_quar_for_tx;
			2'b11 : clk_frm = clk_blf_eigh_for_tx;
		endcase
	end
	else clk_frm = 1'b0;
end


// --- generate clock signal of FM0 Encoder ---
assign clk_fm0 = (m == 2'b00)? clk_blf_for_tx : 1'b0;


// --- generate clock signal of Miller Encoder ---
always@(*) begin
	if(en_tx) begin
		case(m)
			2'b00 : clk_mil = 1'b0;
			2'b01 : clk_mil = clk_blf_for_tx;
			2'b10 : clk_mil = clk_blf_half_for_tx;
			2'b11 : clk_mil = clk_blf_quar_for_tx;
		endcase
	end
	else clk_mil = 1'b0;
end

//----- generate clock signal of Memory -----
always@(negedge clk_frm or negedge rst_n) begin
	if(~rst_n) rd_complete_d <= 1'b0;
	else rd_complete_d <= rd_complete;
end

assign clk_if = clk_frm & en_if & ~rd_complete_d;


endmodule
